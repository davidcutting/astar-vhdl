entity cost is
    port (
        x0, y0 : in std_logic_vector(7 downto 0);
        x, y   : in std_logic_vector(7 downto 0);
        cost   : out std_logic_vector(7 downto 0)
    );
end cost;

architecture Behavioral of cost is

begin

end Behavioral;
